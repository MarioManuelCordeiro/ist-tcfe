.OP 

R1 1 2 1.043096K 
R2 3 2 2.017446K 
R3 2 4 3.136914K 
R4 4 0 4.154300K 
R5 4 5 3.079154K 
R6 0 6 2.025927K 
R7 8 7 1.042267K 
Vo 6 8 0 
H1 4 7 Vo 8.252475K 
G1 5 3 2 4 7.316305m 
Vs 1 0 0.000000 
C 7 5 1.038991u 
.END 
