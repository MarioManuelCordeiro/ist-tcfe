.OP 

R1 1 2 1.015259K 
R2 3 2 2.090689K 
R3 2 4 3.108356K 
R4 4 0 4.101243K 
R5 4 5 3.033480K 
R6 0 6 2.009605K 
R7 8 7 1.005573K 
Vo 6 8 0 
H1 4 7 Vo 8.185741K 
G1 5 3 2 4 7.161103m 
Vs 1 0 0.000000 
Vc 5 7 8.394437 
.END 
